module gnn_accelerator_top_tb();
endmodule
