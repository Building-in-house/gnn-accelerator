module gnn_accelerator_top();
endmodule
